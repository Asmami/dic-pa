    * Pixel sensor
**********************************************************************
**        Copyright (c) 2021 Carsten Wulff Software, Norway
** *******************************************************************
** Created       : wulff at 2021-7-22
** *******************************************************************
**  The MIT License (MIT)
**
**  Permission is hereby granted, free of charge, to any person obtaining a copy
**  of this software and associated documentation files (the "Software"), to deal
**  in the Software without restriction, including without limitation the rights
**  to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
**  copies of the Software, and to permit persons to whom the Software is
**  furnished to do so, subject to the following conditions:
**
**  The above copyright notice and this permission notice shall be included in all
**  copies or substantial portions of the Software.
**
**  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
**  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
**  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
**  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
**  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
**  OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
**  SOFTWARE.
**
**********************************************************************

.SUBCKT PIXEL_SENSOR VBN1 VRAMP VRESET ERASE EXPOSE READ 
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS


XS1 VRESET VSTORE ERASE EXPOSE VDD VSS SENSOR

XC1 VCMP_OUT VSTORE VRAMP VBN1 VDD VSS COMP

XM1 READ VCMP_OUT DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS MEMORY

.ENDS

.SUBCKT MEMORY READ VCMP_OUT
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS

XM1 VCMP_OUT DATA_0 READ VSS MEMCELL
XM2 VCMP_OUT DATA_1 READ VSS MEMCELL
XM3 VCMP_OUT DATA_2 READ VSS MEMCELL
XM4 VCMP_OUT DATA_3 READ VSS MEMCELL
XM5 VCMP_OUT DATA_4 READ VSS MEMCELL
XM6 VCMP_OUT DATA_5 READ VSS MEMCELL
XM7 VCMP_OUT DATA_6 READ VSS MEMCELL
XM8 VCMP_OUT DATA_7 READ VSS MEMCELL

.ENDS

.SUBCKT MEMCELL CMP DATA READ VSS
M1 VG CMP DATA VSS nmos  w=0.2u  l=0.13u
M2 DATA READ DMEM VSS nmos  w=0.4u  l=0.13u
M3 DMEM VG VSS VSS nmos  w=1u  l=0.13u
C1 VG VSS 1p
.ENDS

.SUBCKT SENSOR VRESET VSTORE ERASE EXPOSE VDD VSS
M1 VPG EXPOSE VSTORE VSS nmos w=0.5u l=0.5u
M2 VRESET ERASE VSTORE VSS nmos w=0.5u l=0.5u

* Capacitor to model gate-source capacitance
C1 VSTORE VSS 100f

* Model photocurrent
Rphoto VPG VSS 1G

.ENDS

.SUBCKT COMP VCMP_OUT VSTORE VRAMP VBN1 VDD VSS

* Comparator
M5 VD5 VSTORE VS5 VSS nmos w=0.5u l=0.15u
M6 VS5 VBN1 VSS VSS nmos w=0.5u l=0.5u
M7 VD7 VBN1 VSS VSS nmos w=0.5u l=0.5u
M8 VCMP_OUT VD7 VSS VSS nmos w=0.5u l=0.15u
M9 VD9 VRAMP VS5 VSS nmos w=0.5u l=0.15u

M10 VD9 VD5 VDD VDD pmos w=0.5u l=0.5u
M11 VD5 VD5 VDD VDD pmos w=0.5u l=0.5u
M12 VD7 VD9 VDD VDD pmos w=0.5u l=0.15u
M13 VCMP_OUT VD7 VDD VDD pmos w=0.5u l=0.15u


.ENDS
